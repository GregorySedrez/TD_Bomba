entity bomba is
    port(
		ENTRADA: in bit;
		SAIDA: out bit
    );
end bomba;

architecture arch_bomba of bomba is 
begin
end arch_bomba;